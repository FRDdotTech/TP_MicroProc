LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

entity register_e is
	port (
		CLK, Rin : in std_logic:='0';
		R : in std_logic_vector(8 downto 0);
		Q : out std_logic_vector(8 downto 0):= b"000000000"
	);
end entity;

architecture register_a of register_e is

begin
	
	process (CLK)
	begin
	if rising_edge (CLK) and Rin = '1' then
		Q <= R;
	end if;
	end process;
end architecture;


LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

entity register_bench_e is
end entity;

architecture register_bench_a of register_bench_e is
	component register_e is
		port (
		CLK, Rin : in std_logic:='0';
		R : in std_logic_vector(8 downto 0);
		Q : out std_logic_vector(8 downto 0)
	);
	end component;
	
	signal T_CLK, T_Rin : std_logic:='0';
	signal T_R : std_logic_vector(8 downto 0):= "101010101";
	signal T_Q : std_logic_vector(8 downto 0);
begin
	T_CLK	<= not(T_CLK) after 10 ns;
	T_Rin	<= '1' after 25 ns, '0' after 45 ns, '1' after 65 ns;
	T_R 	<= "000000000" after 47 ns;
	result	: entity work.register_e(register_a) port map(T_CLK, T_Rin, T_R, T_Q);
end architecture;